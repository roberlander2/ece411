import mult_types::*;

module mult_tb;

multiplier_itf itf();

multiplier dut (
    .clk_i          ( itf.clk          ),
    .reset_n_i      ( itf.reset_n      ),
    .multiplicand_i ( itf.multiplicand ),
    .multiplier_i   ( itf.multiplier   ),
    .start_i        ( itf.start        ),
    .ready_o        ( itf.rdy          ),
    .product_o      ( itf.product      ),
    .done_o         ( itf.done         )
);

assign itf.mult_op = dut.ms.op;
default clocking tb_clk @(negedge itf.clk); endclocking

// DO NOT MODIFY CODE ABOVE THIS LINE

/* Uncomment to "monitor" changes to adder operational state over time */
//initial $monitor("dut-op: time: %0t op: %s", $time, dut.ms.op.name);


// Resets the multiplier
task reset();
    itf.reset_n <= 1'b0;
    ##5;
    itf.reset_n <= 1'b1;
    ##1;
endtask : reset

task start();
    itf.start <= 1'b1;
    ##5;
    itf.start <= 1'b0;
    ##1;
endtask : start

// error_e defined in package mult_types in file ../include/types.sv
// Asynchronously reports error in DUT to grading harness
function void report_error(error_e error);
    itf.tb_report_dut_error(error);
endfunction : report_error

initial itf.reset_n = 1'b0;
initial begin
    reset();
    /********************** Your Code Here *****************************/
    //multiply operand
    for (int i = 0; i < 4294967; i++) begin
      for(int j = 0; j < 4294967; j++) begin
        itf.multiplier <= i;
        itf.multiplicand <=j;
        start();
        @(tb_clk iff itf.done == 1'b1);
        assert_equal: assert(itf.product == itf.multiplier * itf.multiplicand)
          else begin
            $error("%0d: %0t: BAD_PRODUCT error detected",`__LINE__,$time);
            report_error(BAD_PRODUCT);
          end
        assert_ready: assert(itf.rdy == 1'b1)
          else begin
            $error("%0d: %0t: NOT_READY error detected",`__LINE__,$time);
            report_error(NOT_READY);
          end
      end
    end

    reset();

    //start and reset coverage while the multiplication is running during the add cycle
    @(tb_clk);
    if(itf.rdy == 1'b1) begin
      start();
    end
    @(tb_clk iff itf.mult_op == ADD);
    start();
    assert(itf.rdy == 1'b0);
    assert(itf.done == 1'b0);
    @(tb_clk iff itf.mult_op == ADD);
    reset();
    assert(itf.rdy == 1'b1)
      else begin
        $error("%0d: %0t: NOT_READY error detected",`__LINE__,$time);
        report_error(NOT_READY);
      end
    assert(itf.done == 1'b0)
      else begin
        $error("%0d: %0t: NOT_READY error detected",`__LINE__,$time);
        report_error(NOT_READY);
      end

      reset();

      //start and reset coverage while the multiplication is running during the shift cycle
      @(tb_clk);
      if(itf.rdy == 1'b1) begin
        start();
      end
      @(tb_clk iff itf.mult_op == SHIFT);
      start();
      assert(itf.rdy == 1'b0);
      assert(itf.done == 1'b0);
      @(tb_clk iff itf.mult_op == SHIFT);
      reset();
      assert(itf.rdy == 1'b1)
        else begin
          $error("%0d: %0t: NOT_READY error detected",`__LINE__,$time);
          report_error(NOT_READY);
        end
      assert(itf.done == 1'b0)
        else begin
          $error("%0d: %0t: NOT_READY error detected",`__LINE__,$time);
          report_error(NOT_READY);
        end



    /*******************************************************************/
    itf.finish(); // Use this finish task in order to let grading harness
                  // complete in process and/or scheduled operations
    $error("Improper Simulation Exit");
end


endmodule : mult_tb
