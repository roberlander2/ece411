module BTB(



);


endmodule: BTB