module mp3(


);

datapath dp

endmodule: mp3