import rv32i_types::*;

module control (
	input clk,
	input rv32i_word inst,
	output control_word_t cw
);


endmodule: control